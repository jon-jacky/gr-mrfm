

//   MRFM Register defines

`define FR_MRFM_DECIM             7'd64
`define FR_MRFM_FREQ              7'd65
`define FR_MRFM_PHASE             7'd66
`define FR_MRFM_IIR_COEFF         7'd67
`define FR_MRFM_IIR_SHIFT         7'd68
`define FR_MRFM_DEBUG             7'd69
`define FR_MRFM_COMP_A11          7'd70
`define FR_MRFM_COMP_A12          7'd71
`define FR_MRFM_COMP_A21          7'd72
`define FR_MRFM_COMP_A22          7'd73
`define FR_MRFM_COMP_SHIFT        7'd74
`define FR_MRFM_SCALE_K0          7'd75
`define FR_MRFM_SCALE_K1          7'd76
`define FR_USER_13                7'd77
`define FR_USER_14                7'd78
`define FR_USER_15                7'd79

